
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017
signal mem : ram_t := (

--			***** COLOR PALLETE *****


	
		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00D4BC00", -- R: 0 G: 188 B: 212
		2 =>	x"001E6933", -- R: 51 G: 105 B: 30
		3 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		4 =>	x"004AC38B", -- R: 139 G: 195 B: 74
		5 =>	x"00205E1B", -- R: 27 G: 94 B: 32
		6 =>	x"000C66A6", -- R: 166 G: 102 B: 12
		7 =>	x"00152A38", -- R: 56 G: 42 B: 21
		8 =>	x"000A0A0A", -- R: 10 G: 10 B: 10
		9 =>	x"001A1A1A", -- R: 26 G: 26 B: 26
		10 =>	x"000B0B0B", -- R: 11 G: 11 B: 11
		11 =>	x"0092CD90", -- R: 144 G: 205 B: 146
		12 =>	x"0050AF4C", -- R: 76 G: 175 B: 80
		13 =>	x"0066B963", -- R: 99 G: 185 B: 102
		14 =>	x"002257FF", -- R: 255 G: 87 B: 34
		15 =>	x"000098FF", -- R: 255 G: 152 B: 0
		16 =>	x"00D7BC07", -- R: 7 G: 188 B: 215
		17 =>	x"00020202", -- R: 2 G: 2 B: 2
		18 =>	x"00010101", -- R: 1 G: 1 B: 1
		19 =>	x"00000000", -- Unused
		20 =>	x"00000000", -- Unused
		21 =>	x"00000000", -- Unused
		22 =>	x"00000000", -- Unused
		23 =>	x"00000000", -- Unused
		24 =>	x"00000000", -- Unused
		25 =>	x"00000000", -- Unused
		26 =>	x"00000000", -- Unused
		27 =>	x"00000000", -- Unused
		28 =>	x"00000000", -- Unused
		29 =>	x"00000000", -- Unused
		30 =>	x"00000000", -- Unused
		31 =>	x"00000000", -- Unused
		32 =>	x"00000000", -- Unused
		33 =>	x"00000000", -- Unused
		34 =>	x"00000000", -- Unused
		35 =>	x"00000000", -- Unused
		36 =>	x"00000000", -- Unused
		37 =>	x"00000000", -- Unused
		38 =>	x"00000000", -- Unused
		39 =>	x"00000000", -- Unused
		40 =>	x"00000000", -- Unused
		41 =>	x"00000000", -- Unused
		42 =>	x"00000000", -- Unused
		43 =>	x"00000000", -- Unused
		44 =>	x"00000000", -- Unused
		45 =>	x"00000000", -- Unused
		46 =>	x"00000000", -- Unused
		47 =>	x"00000000", -- Unused
		48 =>	x"00000000", -- Unused
		49 =>	x"00000000", -- Unused
		50 =>	x"00000000", -- Unused
		51 =>	x"00000000", -- Unused
		52 =>	x"00000000", -- Unused
		53 =>	x"00000000", -- Unused
		54 =>	x"00000000", -- Unused
		55 =>	x"00000000", -- Unused
		56 =>	x"00000000", -- Unused
		57 =>	x"00000000", -- Unused
		58 =>	x"00000000", -- Unused
		59 =>	x"00000000", -- Unused
		60 =>	x"00000000", -- Unused
		61 =>	x"00000000", -- Unused
		62 =>	x"00000000", -- Unused
		63 =>	x"00000000", -- Unused
		64 =>	x"00000000", -- Unused
		65 =>	x"00000000", -- Unused
		66 =>	x"00000000", -- Unused
		67 =>	x"00000000", -- Unused
		68 =>	x"00000000", -- Unused
		69 =>	x"00000000", -- Unused
		70 =>	x"00000000", -- Unused
		71 =>	x"00000000", -- Unused
		72 =>	x"00000000", -- Unused
		73 =>	x"00000000", -- Unused
		74 =>	x"00000000", -- Unused
		75 =>	x"00000000", -- Unused
		76 =>	x"00000000", -- Unused
		77 =>	x"00000000", -- Unused
		78 =>	x"00000000", -- Unused
		79 =>	x"00000000", -- Unused
		80 =>	x"00000000", -- Unused
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused


		
--			***** 16x16 IMAGES *****
		
		
				255 =>	x"01010101", -- IMG_16x16_bg00
		256 =>	x"01010101",
		257 =>	x"01010101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01010101",
		261 =>	x"01010101",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01010101",
		265 =>	x"01010101",
		266 =>	x"01010101",
		267 =>	x"01010101",
		268 =>	x"01010101",
		269 =>	x"01010101",
		270 =>	x"01010101",
		271 =>	x"01010101",
		272 =>	x"01020101",
		273 =>	x"01010101",
		274 =>	x"02020101",
		275 =>	x"01010101",
		276 =>	x"01020101",
		277 =>	x"01010101",
		278 =>	x"02020201",
		279 =>	x"01010101",
		280 =>	x"02020203",
		281 =>	x"03010101",
		282 =>	x"01020202",
		283 =>	x"01010101",
		284 =>	x"02040203",
		285 =>	x"03030101",
		286 =>	x"01020202",
		287 =>	x"01010101",
		288 =>	x"02040202",
		289 =>	x"03030303",
		290 =>	x"01010204",
		291 =>	x"01010202",
		292 =>	x"04040402",
		293 =>	x"02030303",
		294 =>	x"01010204",
		295 =>	x"04020204",
		296 =>	x"04040404",
		297 =>	x"02020303",
		298 =>	x"01010204",
		299 =>	x"02020404",
		300 =>	x"04040404",
		301 =>	x"04040203",
		302 =>	x"03010204",
		303 =>	x"02040404",
		304 =>	x"04040404",
		305 =>	x"04040402",
		306 =>	x"03010204",
		307 =>	x"04040404",
		308 =>	x"04040404",
		309 =>	x"04040402",
		310 =>	x"04020204",
		311 =>	x"04040404",
		312 =>	x"04040404",
		313 =>	x"04040404",
		314 =>	x"04040404",
		315 =>	x"04040404",
		316 =>	x"04040404",
		317 =>	x"04040404",
		318 =>	x"04040404",
		319 =>	x"01010101", -- IMG_16x16_bg01
		320 =>	x"01010101",
		321 =>	x"01010101",
		322 =>	x"01010101",
		323 =>	x"01010101",
		324 =>	x"01010101",
		325 =>	x"01010101",
		326 =>	x"01010101",
		327 =>	x"01010101",
		328 =>	x"01010101",
		329 =>	x"01010101",
		330 =>	x"01010101",
		331 =>	x"01010101",
		332 =>	x"01010101",
		333 =>	x"01010101",
		334 =>	x"01010101",
		335 =>	x"01010101",
		336 =>	x"01010101",
		337 =>	x"01010101",
		338 =>	x"01020201",
		339 =>	x"03010101",
		340 =>	x"01010101",
		341 =>	x"01010101",
		342 =>	x"02020101",
		343 =>	x"03030101",
		344 =>	x"01010101",
		345 =>	x"01010102",
		346 =>	x"02030101",
		347 =>	x"02030301",
		348 =>	x"01010101",
		349 =>	x"01010204",
		350 =>	x"02030101",
		351 =>	x"02030303",
		352 =>	x"01010101",
		353 =>	x"01020402",
		354 =>	x"02030101",
		355 =>	x"04020303",
		356 =>	x"03010101",
		357 =>	x"01020402",
		358 =>	x"03030101",
		359 =>	x"04040303",
		360 =>	x"03010101",
		361 =>	x"01040404",
		362 =>	x"02030301",
		363 =>	x"04040203",
		364 =>	x"03030402",
		365 =>	x"04040404",
		366 =>	x"02040301",
		367 =>	x"04040202",
		368 =>	x"03030402",
		369 =>	x"04040404",
		370 =>	x"04040101",
		371 =>	x"04040404",
		372 =>	x"04040404",
		373 =>	x"04040404",
		374 =>	x"04040404",
		375 =>	x"04040404",
		376 =>	x"04040404",
		377 =>	x"04040404",
		378 =>	x"04040404",
		379 =>	x"04040404",
		380 =>	x"04040404",
		381 =>	x"04040404",
		382 =>	x"04040404",
		383 =>	x"01010101", -- IMG_16x16_bg02
		384 =>	x"01010101",
		385 =>	x"01010101",
		386 =>	x"01010101",
		387 =>	x"01010101",
		388 =>	x"01010101",
		389 =>	x"01010101",
		390 =>	x"01010101",
		391 =>	x"01010101",
		392 =>	x"01020101",
		393 =>	x"01010101",
		394 =>	x"01010101",
		395 =>	x"01010101",
		396 =>	x"02020101",
		397 =>	x"01010101",
		398 =>	x"01010102",
		399 =>	x"01010101",
		400 =>	x"02020101",
		401 =>	x"01010101",
		402 =>	x"01010102",
		403 =>	x"01010101",
		404 =>	x"02020101",
		405 =>	x"01010101",
		406 =>	x"01010101",
		407 =>	x"01010101",
		408 =>	x"02020201",
		409 =>	x"01010101",
		410 =>	x"01010101",
		411 =>	x"01010101",
		412 =>	x"02040203",
		413 =>	x"01010101",
		414 =>	x"01010102",
		415 =>	x"01010101",
		416 =>	x"02040203",
		417 =>	x"03010101",
		418 =>	x"01010102",
		419 =>	x"01010101",
		420 =>	x"02040203",
		421 =>	x"03010101",
		422 =>	x"01010102",
		423 =>	x"01010102",
		424 =>	x"02040402",
		425 =>	x"03030101",
		426 =>	x"01010102",
		427 =>	x"01040202",
		428 =>	x"04040402",
		429 =>	x"02040303",
		430 =>	x"01010204",
		431 =>	x"01040404",
		432 =>	x"04040404",
		433 =>	x"02020403",
		434 =>	x"01020404",
		435 =>	x"04040404",
		436 =>	x"04040404",
		437 =>	x"04020204",
		438 =>	x"01020404",
		439 =>	x"04040404",
		440 =>	x"04040404",
		441 =>	x"04040404",
		442 =>	x"04040404",
		443 =>	x"04040404",
		444 =>	x"04040404",
		445 =>	x"04040404",
		446 =>	x"04040404",
		447 =>	x"04040404", -- IMG_16x16_bg10
		448 =>	x"04040404",
		449 =>	x"04040404",
		450 =>	x"04040404",
		451 =>	x"04040404",
		452 =>	x"04040404",
		453 =>	x"04040404",
		454 =>	x"04040404",
		455 =>	x"04040404",
		456 =>	x"04040404",
		457 =>	x"04040404",
		458 =>	x"04040404",
		459 =>	x"04040404",
		460 =>	x"04040404",
		461 =>	x"04040404",
		462 =>	x"04040404",
		463 =>	x"04040404",
		464 =>	x"04040404",
		465 =>	x"04040404",
		466 =>	x"04040404",
		467 =>	x"04040404",
		468 =>	x"04040404",
		469 =>	x"04040404",
		470 =>	x"04040404",
		471 =>	x"04040404",
		472 =>	x"04040404",
		473 =>	x"04040404",
		474 =>	x"04040404",
		475 =>	x"04040404",
		476 =>	x"04040404",
		477 =>	x"04040404",
		478 =>	x"04040404",
		479 =>	x"04040404",
		480 =>	x"04040404",
		481 =>	x"04040404",
		482 =>	x"04040404",
		483 =>	x"04040404",
		484 =>	x"04040404",
		485 =>	x"04040404",
		486 =>	x"04040404",
		487 =>	x"04040404",
		488 =>	x"04040404",
		489 =>	x"04040404",
		490 =>	x"04040404",
		491 =>	x"04040404",
		492 =>	x"04040404",
		493 =>	x"04040404",
		494 =>	x"04040404",
		495 =>	x"04040404",
		496 =>	x"04040404",
		497 =>	x"04040404",
		498 =>	x"04040404",
		499 =>	x"04040404",
		500 =>	x"04040404",
		501 =>	x"04040404",
		502 =>	x"04040404",
		503 =>	x"04040404",
		504 =>	x"04040404",
		505 =>	x"04040404",
		506 =>	x"04040404",
		507 =>	x"04040404",
		508 =>	x"04040404",
		509 =>	x"04040404",
		510 =>	x"04040404",
		511 =>	x"04040404", -- IMG_16x16_bg11
		512 =>	x"04040404",
		513 =>	x"04040404",
		514 =>	x"04040404",
		515 =>	x"04040404",
		516 =>	x"04040404",
		517 =>	x"04040404",
		518 =>	x"04040404",
		519 =>	x"04040404",
		520 =>	x"04040404",
		521 =>	x"04040404",
		522 =>	x"04040404",
		523 =>	x"04040404",
		524 =>	x"04040404",
		525 =>	x"04040504",
		526 =>	x"04040404",
		527 =>	x"04040404",
		528 =>	x"04040404",
		529 =>	x"04040505",
		530 =>	x"04040404",
		531 =>	x"04040404",
		532 =>	x"04040404",
		533 =>	x"04040405",
		534 =>	x"04040404",
		535 =>	x"04040404",
		536 =>	x"04040404",
		537 =>	x"04040405",
		538 =>	x"04040404",
		539 =>	x"04040404",
		540 =>	x"04040404",
		541 =>	x"04040405",
		542 =>	x"04040404",
		543 =>	x"04040404",
		544 =>	x"04040404",
		545 =>	x"04040405",
		546 =>	x"04040404",
		547 =>	x"04040404",
		548 =>	x"04040404",
		549 =>	x"04040505",
		550 =>	x"04040404",
		551 =>	x"04040404",
		552 =>	x"04040404",
		553 =>	x"04040505",
		554 =>	x"04040404",
		555 =>	x"04040404",
		556 =>	x"04040404",
		557 =>	x"04050504",
		558 =>	x"04040404",
		559 =>	x"04040404",
		560 =>	x"04040404",
		561 =>	x"05050404",
		562 =>	x"04040404",
		563 =>	x"04040404",
		564 =>	x"04040404",
		565 =>	x"05050404",
		566 =>	x"04040404",
		567 =>	x"04040404",
		568 =>	x"04040405",
		569 =>	x"05050404",
		570 =>	x"04040404",
		571 =>	x"04040404",
		572 =>	x"04040405",
		573 =>	x"05040404",
		574 =>	x"04040404",
		575 =>	x"04040404", -- IMG_16x16_bg12
		576 =>	x"04040404",
		577 =>	x"04040404",
		578 =>	x"04040404",
		579 =>	x"04040404",
		580 =>	x"04040404",
		581 =>	x"04040404",
		582 =>	x"04040404",
		583 =>	x"04040404",
		584 =>	x"04040404",
		585 =>	x"04040404",
		586 =>	x"04040404",
		587 =>	x"04040404",
		588 =>	x"04040404",
		589 =>	x"04040505",
		590 =>	x"04040404",
		591 =>	x"04040404",
		592 =>	x"04040404",
		593 =>	x"04040405",
		594 =>	x"04040404",
		595 =>	x"04040404",
		596 =>	x"04040404",
		597 =>	x"04040405",
		598 =>	x"04040404",
		599 =>	x"04040404",
		600 =>	x"04040404",
		601 =>	x"04040505",
		602 =>	x"04040404",
		603 =>	x"04040404",
		604 =>	x"04040404",
		605 =>	x"04040505",
		606 =>	x"04040404",
		607 =>	x"04040404",
		608 =>	x"04040404",
		609 =>	x"04040505",
		610 =>	x"04040404",
		611 =>	x"04040404",
		612 =>	x"04040404",
		613 =>	x"04040505",
		614 =>	x"05040404",
		615 =>	x"04040404",
		616 =>	x"04040404",
		617 =>	x"04040405",
		618 =>	x"05040404",
		619 =>	x"04040404",
		620 =>	x"04040404",
		621 =>	x"04040405",
		622 =>	x"05050404",
		623 =>	x"04040404",
		624 =>	x"04040404",
		625 =>	x"04040405",
		626 =>	x"05050404",
		627 =>	x"04040404",
		628 =>	x"04040404",
		629 =>	x"04040404",
		630 =>	x"05050504",
		631 =>	x"04040404",
		632 =>	x"04040404",
		633 =>	x"04040404",
		634 =>	x"04050504",
		635 =>	x"04040404",
		636 =>	x"04040404",
		637 =>	x"04040404",
		638 =>	x"04050404",
		639 =>	x"04040404", -- IMG_16x16_bg20
		640 =>	x"04040404",
		641 =>	x"04040404",
		642 =>	x"04040404",
		643 =>	x"04040404",
		644 =>	x"04040404",
		645 =>	x"04040404",
		646 =>	x"04040404",
		647 =>	x"04040404",
		648 =>	x"04040404",
		649 =>	x"04040404",
		650 =>	x"04040404",
		651 =>	x"04040404",
		652 =>	x"04040404",
		653 =>	x"04040404",
		654 =>	x"04040404",
		655 =>	x"04040404",
		656 =>	x"04040404",
		657 =>	x"04040404",
		658 =>	x"04040404",
		659 =>	x"04040404",
		660 =>	x"04040404",
		661 =>	x"04040404",
		662 =>	x"04040404",
		663 =>	x"04040404",
		664 =>	x"04040404",
		665 =>	x"04040404",
		666 =>	x"04040404",
		667 =>	x"04040404",
		668 =>	x"04040404",
		669 =>	x"04040404",
		670 =>	x"04040404",
		671 =>	x"04040404",
		672 =>	x"04040404",
		673 =>	x"04040404",
		674 =>	x"04040404",
		675 =>	x"04040404",
		676 =>	x"04040404",
		677 =>	x"04040404",
		678 =>	x"04040404",
		679 =>	x"04040404",
		680 =>	x"04040404",
		681 =>	x"04040404",
		682 =>	x"04040404",
		683 =>	x"04040404",
		684 =>	x"04040404",
		685 =>	x"04040404",
		686 =>	x"04040404",
		687 =>	x"04040404",
		688 =>	x"04040404",
		689 =>	x"04040404",
		690 =>	x"04040404",
		691 =>	x"04040404",
		692 =>	x"04040404",
		693 =>	x"04040205",
		694 =>	x"04040404",
		695 =>	x"04040404",
		696 =>	x"04040404",
		697 =>	x"04040405",
		698 =>	x"04040404",
		699 =>	x"04040404",
		700 =>	x"04040404",
		701 =>	x"04040205",
		702 =>	x"04040404",
		703 =>	x"04040404", -- IMG_16x16_bg21
		704 =>	x"04040405",
		705 =>	x"05040404",
		706 =>	x"04040404",
		707 =>	x"04040404",
		708 =>	x"04040405",
		709 =>	x"05040404",
		710 =>	x"04040404",
		711 =>	x"04040404",
		712 =>	x"04040405",
		713 =>	x"05040404",
		714 =>	x"04040404",
		715 =>	x"04040404",
		716 =>	x"04040404",
		717 =>	x"05040404",
		718 =>	x"04040404",
		719 =>	x"04040404",
		720 =>	x"04040405",
		721 =>	x"05040404",
		722 =>	x"04040404",
		723 =>	x"04040404",
		724 =>	x"04040405",
		725 =>	x"04040404",
		726 =>	x"04040404",
		727 =>	x"04040404",
		728 =>	x"04040404",
		729 =>	x"04040404",
		730 =>	x"04040404",
		731 =>	x"04040404",
		732 =>	x"04040404",
		733 =>	x"04040404",
		734 =>	x"04040404",
		735 =>	x"04040404",
		736 =>	x"04040404",
		737 =>	x"04040404",
		738 =>	x"04040404",
		739 =>	x"04040404",
		740 =>	x"04040404",
		741 =>	x"04040404",
		742 =>	x"04040404",
		743 =>	x"04040404",
		744 =>	x"04040404",
		745 =>	x"04040404",
		746 =>	x"04040404",
		747 =>	x"04040404",
		748 =>	x"04040404",
		749 =>	x"04040404",
		750 =>	x"04040404",
		751 =>	x"04040404",
		752 =>	x"04040404",
		753 =>	x"04040404",
		754 =>	x"04040404",
		755 =>	x"04040404",
		756 =>	x"04040404",
		757 =>	x"04040404",
		758 =>	x"04040404",
		759 =>	x"04040404",
		760 =>	x"04040404",
		761 =>	x"04040404",
		762 =>	x"04040404",
		763 =>	x"04040404",
		764 =>	x"04040404",
		765 =>	x"04040404",
		766 =>	x"04040404",
		767 =>	x"04040404", -- IMG_16x16_bg22
		768 =>	x"04040404",
		769 =>	x"04040404",
		770 =>	x"04050404",
		771 =>	x"04040404",
		772 =>	x"04040404",
		773 =>	x"04040404",
		774 =>	x"05050404",
		775 =>	x"04040404",
		776 =>	x"04040404",
		777 =>	x"04040404",
		778 =>	x"05050404",
		779 =>	x"04040404",
		780 =>	x"04040404",
		781 =>	x"04040404",
		782 =>	x"04040404",
		783 =>	x"04040404",
		784 =>	x"04040404",
		785 =>	x"04040404",
		786 =>	x"04040404",
		787 =>	x"04040404",
		788 =>	x"04040404",
		789 =>	x"04040404",
		790 =>	x"04040404",
		791 =>	x"04040404",
		792 =>	x"04040404",
		793 =>	x"04040404",
		794 =>	x"04040404",
		795 =>	x"04040404",
		796 =>	x"04040404",
		797 =>	x"04040404",
		798 =>	x"04040404",
		799 =>	x"04040404",
		800 =>	x"04040404",
		801 =>	x"04040404",
		802 =>	x"04040404",
		803 =>	x"04040404",
		804 =>	x"04040404",
		805 =>	x"04040404",
		806 =>	x"04040404",
		807 =>	x"04040404",
		808 =>	x"04040404",
		809 =>	x"04040404",
		810 =>	x"04040404",
		811 =>	x"04040404",
		812 =>	x"04040404",
		813 =>	x"04040404",
		814 =>	x"04040404",
		815 =>	x"04040404",
		816 =>	x"04040404",
		817 =>	x"04040404",
		818 =>	x"04040404",
		819 =>	x"04040404",
		820 =>	x"04040404",
		821 =>	x"04040404",
		822 =>	x"04040404",
		823 =>	x"05050404",
		824 =>	x"04040404",
		825 =>	x"04040404",
		826 =>	x"04040404",
		827 =>	x"04050204",
		828 =>	x"04040404",
		829 =>	x"04040404",
		830 =>	x"04040404",
		831 =>	x"04040404", -- IMG_16x16_bg30
		832 =>	x"04040404",
		833 =>	x"04020504",
		834 =>	x"04040404",
		835 =>	x"04040404",
		836 =>	x"04040404",
		837 =>	x"04040504",
		838 =>	x"04040404",
		839 =>	x"04040404",
		840 =>	x"04040404",
		841 =>	x"04020504",
		842 =>	x"04040404",
		843 =>	x"04040404",
		844 =>	x"04040404",
		845 =>	x"02050504",
		846 =>	x"04040404",
		847 =>	x"04040404",
		848 =>	x"04040404",
		849 =>	x"05020404",
		850 =>	x"04040404",
		851 =>	x"04040404",
		852 =>	x"04040405",
		853 =>	x"05040404",
		854 =>	x"04040404",
		855 =>	x"04040404",
		856 =>	x"04040405",
		857 =>	x"02040404",
		858 =>	x"04040404",
		859 =>	x"04040404",
		860 =>	x"04040405",
		861 =>	x"02040404",
		862 =>	x"04040404",
		863 =>	x"04040404",
		864 =>	x"04040504",
		865 =>	x"04040404",
		866 =>	x"04040404",
		867 =>	x"04040404",
		868 =>	x"04050504",
		869 =>	x"04040404",
		870 =>	x"04040404",
		871 =>	x"04040404",
		872 =>	x"04050204",
		873 =>	x"04040404",
		874 =>	x"04040404",
		875 =>	x"04040404",
		876 =>	x"04050204",
		877 =>	x"04040404",
		878 =>	x"04040404",
		879 =>	x"04040404",
		880 =>	x"05050404",
		881 =>	x"04040404",
		882 =>	x"04040404",
		883 =>	x"04040404",
		884 =>	x"04040404",
		885 =>	x"04040404",
		886 =>	x"04040404",
		887 =>	x"04040404",
		888 =>	x"04040404",
		889 =>	x"04040404",
		890 =>	x"04040404",
		891 =>	x"04040404",
		892 =>	x"04040404",
		893 =>	x"04040404",
		894 =>	x"04040404",
		895 =>	x"04040404", -- IMG_16x16_bg31
		896 =>	x"04040404",
		897 =>	x"04040404",
		898 =>	x"04040404",
		899 =>	x"04040404",
		900 =>	x"04040404",
		901 =>	x"04040404",
		902 =>	x"04040404",
		903 =>	x"04040404",
		904 =>	x"04040404",
		905 =>	x"04040404",
		906 =>	x"04040404",
		907 =>	x"04040404",
		908 =>	x"04040404",
		909 =>	x"04040404",
		910 =>	x"04040404",
		911 =>	x"04040404",
		912 =>	x"04040404",
		913 =>	x"04040404",
		914 =>	x"04040404",
		915 =>	x"04040404",
		916 =>	x"04040404",
		917 =>	x"04040404",
		918 =>	x"04040404",
		919 =>	x"04040404",
		920 =>	x"04040404",
		921 =>	x"04040404",
		922 =>	x"04040404",
		923 =>	x"04040404",
		924 =>	x"04040404",
		925 =>	x"04040404",
		926 =>	x"04040404",
		927 =>	x"04040404",
		928 =>	x"04040404",
		929 =>	x"04040404",
		930 =>	x"04040404",
		931 =>	x"04040404",
		932 =>	x"04040404",
		933 =>	x"04040404",
		934 =>	x"04040404",
		935 =>	x"04040404",
		936 =>	x"04040404",
		937 =>	x"04040404",
		938 =>	x"04040404",
		939 =>	x"04040404",
		940 =>	x"04040404",
		941 =>	x"04040404",
		942 =>	x"04040404",
		943 =>	x"04040404",
		944 =>	x"04040404",
		945 =>	x"04040404",
		946 =>	x"04040404",
		947 =>	x"04040404",
		948 =>	x"04040404",
		949 =>	x"04040404",
		950 =>	x"04040404",
		951 =>	x"04040404",
		952 =>	x"04040404",
		953 =>	x"04040404",
		954 =>	x"04040404",
		955 =>	x"04040404",
		956 =>	x"04040404",
		957 =>	x"04040404",
		958 =>	x"04040404",
		959 =>	x"04050204", -- IMG_16x16_bg32
		960 =>	x"04040404",
		961 =>	x"04040404",
		962 =>	x"04040404",
		963 =>	x"02050204",
		964 =>	x"04040404",
		965 =>	x"04040404",
		966 =>	x"04040404",
		967 =>	x"04050204",
		968 =>	x"04040404",
		969 =>	x"04040404",
		970 =>	x"04040404",
		971 =>	x"04050204",
		972 =>	x"04040404",
		973 =>	x"04040404",
		974 =>	x"04040404",
		975 =>	x"04050204",
		976 =>	x"04040404",
		977 =>	x"04040404",
		978 =>	x"04040404",
		979 =>	x"04050504",
		980 =>	x"04040404",
		981 =>	x"04040404",
		982 =>	x"04040404",
		983 =>	x"04040504",
		984 =>	x"04040404",
		985 =>	x"04040404",
		986 =>	x"04040404",
		987 =>	x"04040505",
		988 =>	x"04040404",
		989 =>	x"04040404",
		990 =>	x"04040404",
		991 =>	x"04040205",
		992 =>	x"04040404",
		993 =>	x"04040404",
		994 =>	x"04040404",
		995 =>	x"04040405",
		996 =>	x"05040404",
		997 =>	x"04040404",
		998 =>	x"04040404",
		999 =>	x"04040404",
		1000 =>	x"05040404",
		1001 =>	x"04040404",
		1002 =>	x"04040404",
		1003 =>	x"04040404",
		1004 =>	x"05050404",
		1005 =>	x"04040404",
		1006 =>	x"04040404",
		1007 =>	x"04040404",
		1008 =>	x"02050404",
		1009 =>	x"04040404",
		1010 =>	x"04040404",
		1011 =>	x"04040404",
		1012 =>	x"04050404",
		1013 =>	x"04040404",
		1014 =>	x"04040404",
		1015 =>	x"04040404",
		1016 =>	x"04050404",
		1017 =>	x"04040404",
		1018 =>	x"04040404",
		1019 =>	x"04040404",
		1020 =>	x"04050404",
		1021 =>	x"04040404",
		1022 =>	x"04040404",
		1023 =>	x"04040404", -- IMG_16x16_bg40
		1024 =>	x"04040404",
		1025 =>	x"04040404",
		1026 =>	x"04040404",
		1027 =>	x"04040404",
		1028 =>	x"04040404",
		1029 =>	x"04040404",
		1030 =>	x"04040404",
		1031 =>	x"04040404",
		1032 =>	x"04040404",
		1033 =>	x"04040404",
		1034 =>	x"04040404",
		1035 =>	x"04040404",
		1036 =>	x"04040404",
		1037 =>	x"04040404",
		1038 =>	x"04040404",
		1039 =>	x"04040404",
		1040 =>	x"04040404",
		1041 =>	x"04040404",
		1042 =>	x"04040404",
		1043 =>	x"04040404",
		1044 =>	x"04040404",
		1045 =>	x"04040404",
		1046 =>	x"04040404",
		1047 =>	x"04040404",
		1048 =>	x"04040404",
		1049 =>	x"04040404",
		1050 =>	x"04040404",
		1051 =>	x"04040404",
		1052 =>	x"04040404",
		1053 =>	x"04040404",
		1054 =>	x"04040404",
		1055 =>	x"04040404",
		1056 =>	x"04040400",
		1057 =>	x"00040404",
		1058 =>	x"04040404",
		1059 =>	x"04040404",
		1060 =>	x"00000000",
		1061 =>	x"00000000",
		1062 =>	x"04040404",
		1063 =>	x"00000000",
		1064 =>	x"00000606",
		1065 =>	x"06060600",
		1066 =>	x"00000000",
		1067 =>	x"06060606",
		1068 =>	x"06060606",
		1069 =>	x"06060606",
		1070 =>	x"06060606",
		1071 =>	x"06060606",
		1072 =>	x"06060606",
		1073 =>	x"06060606",
		1074 =>	x"06060606",
		1075 =>	x"06060606",
		1076 =>	x"06060606",
		1077 =>	x"06060606",
		1078 =>	x"06060606",
		1079 =>	x"06060606",
		1080 =>	x"06060606",
		1081 =>	x"06060606",
		1082 =>	x"06060606",
		1083 =>	x"06060606",
		1084 =>	x"06060606",
		1085 =>	x"06060606",
		1086 =>	x"06060606",
		1087 =>	x"04040404", -- IMG_16x16_bg41
		1088 =>	x"04040404",
		1089 =>	x"04040404",
		1090 =>	x"04040404",
		1091 =>	x"04040404",
		1092 =>	x"04040404",
		1093 =>	x"04040404",
		1094 =>	x"04040404",
		1095 =>	x"04040404",
		1096 =>	x"04040404",
		1097 =>	x"04040404",
		1098 =>	x"04040404",
		1099 =>	x"04040404",
		1100 =>	x"04040404",
		1101 =>	x"04040404",
		1102 =>	x"04040404",
		1103 =>	x"04040404",
		1104 =>	x"04040404",
		1105 =>	x"04040404",
		1106 =>	x"04040404",
		1107 =>	x"04040404",
		1108 =>	x"04040404",
		1109 =>	x"04040404",
		1110 =>	x"04040404",
		1111 =>	x"04040404",
		1112 =>	x"04040404",
		1113 =>	x"04040404",
		1114 =>	x"04040404",
		1115 =>	x"04040404",
		1116 =>	x"04040404",
		1117 =>	x"04040404",
		1118 =>	x"04040404",
		1119 =>	x"04040404",
		1120 =>	x"04040404",
		1121 =>	x"00040404",
		1122 =>	x"04040404",
		1123 =>	x"04040404",
		1124 =>	x"04000000",
		1125 =>	x"00000004",
		1126 =>	x"04040404",
		1127 =>	x"00000000",
		1128 =>	x"00060606",
		1129 =>	x"06060600",
		1130 =>	x"00000000",
		1131 =>	x"06060606",
		1132 =>	x"06060606",
		1133 =>	x"06060606",
		1134 =>	x"06060606",
		1135 =>	x"06060606",
		1136 =>	x"06060606",
		1137 =>	x"06060606",
		1138 =>	x"06060606",
		1139 =>	x"06060606",
		1140 =>	x"06060606",
		1141 =>	x"06060606",
		1142 =>	x"06060606",
		1143 =>	x"06060606",
		1144 =>	x"06060606",
		1145 =>	x"06060606",
		1146 =>	x"06060606",
		1147 =>	x"06060606",
		1148 =>	x"06060606",
		1149 =>	x"06060606",
		1150 =>	x"06060606",
		1151 =>	x"04040404", -- IMG_16x16_bg42
		1152 =>	x"04050404",
		1153 =>	x"04040404",
		1154 =>	x"04040404",
		1155 =>	x"04040404",
		1156 =>	x"04040404",
		1157 =>	x"04040404",
		1158 =>	x"04040404",
		1159 =>	x"04040404",
		1160 =>	x"04040404",
		1161 =>	x"04040404",
		1162 =>	x"04040404",
		1163 =>	x"04040404",
		1164 =>	x"04040404",
		1165 =>	x"04040404",
		1166 =>	x"04040404",
		1167 =>	x"04040404",
		1168 =>	x"04040404",
		1169 =>	x"04040404",
		1170 =>	x"04040404",
		1171 =>	x"04040404",
		1172 =>	x"04040404",
		1173 =>	x"04040404",
		1174 =>	x"04040404",
		1175 =>	x"04040404",
		1176 =>	x"04040404",
		1177 =>	x"04040404",
		1178 =>	x"04040404",
		1179 =>	x"04040404",
		1180 =>	x"04040404",
		1181 =>	x"04040404",
		1182 =>	x"04040404",
		1183 =>	x"04040404",
		1184 =>	x"00000004",
		1185 =>	x"04040404",
		1186 =>	x"04040404",
		1187 =>	x"00000000",
		1188 =>	x"00000000",
		1189 =>	x"00040404",
		1190 =>	x"04040404",
		1191 =>	x"00060606",
		1192 =>	x"06060606",
		1193 =>	x"00000000",
		1194 =>	x"00000000",
		1195 =>	x"06060606",
		1196 =>	x"06060606",
		1197 =>	x"06060606",
		1198 =>	x"06000006",
		1199 =>	x"06060606",
		1200 =>	x"06060606",
		1201 =>	x"06060606",
		1202 =>	x"06060606",
		1203 =>	x"06060606",
		1204 =>	x"06060606",
		1205 =>	x"06060606",
		1206 =>	x"06060606",
		1207 =>	x"06060606",
		1208 =>	x"06060606",
		1209 =>	x"06060606",
		1210 =>	x"06060606",
		1211 =>	x"06060606",
		1212 =>	x"06060606",
		1213 =>	x"06060606",
		1214 =>	x"06060606",
		1215 =>	x"06060606", -- IMG_16x16_bg50
		1216 =>	x"06060606",
		1217 =>	x"06060606",
		1218 =>	x"06060606",
		1219 =>	x"06060606",
		1220 =>	x"06060606",
		1221 =>	x"06060606",
		1222 =>	x"06060606",
		1223 =>	x"06060606",
		1224 =>	x"06060606",
		1225 =>	x"06060606",
		1226 =>	x"06060606",
		1227 =>	x"06060606",
		1228 =>	x"06060606",
		1229 =>	x"06060606",
		1230 =>	x"06060606",
		1231 =>	x"06060606",
		1232 =>	x"06060606",
		1233 =>	x"06060606",
		1234 =>	x"07070606",
		1235 =>	x"06060606",
		1236 =>	x"06060606",
		1237 =>	x"06060606",
		1238 =>	x"06070707",
		1239 =>	x"06060606",
		1240 =>	x"06060606",
		1241 =>	x"06060606",
		1242 =>	x"06060606",
		1243 =>	x"06060606",
		1244 =>	x"06060606",
		1245 =>	x"06060606",
		1246 =>	x"06060606",
		1247 =>	x"06060606",
		1248 =>	x"06060606",
		1249 =>	x"06060606",
		1250 =>	x"06060607",
		1251 =>	x"06060606",
		1252 =>	x"06060606",
		1253 =>	x"06060606",
		1254 =>	x"06060606",
		1255 =>	x"06060606",
		1256 =>	x"06060606",
		1257 =>	x"06060606",
		1258 =>	x"06060606",
		1259 =>	x"06060606",
		1260 =>	x"06060606",
		1261 =>	x"06060606",
		1262 =>	x"06060606",
		1263 =>	x"06060606",
		1264 =>	x"06060606",
		1265 =>	x"06060606",
		1266 =>	x"06060606",
		1267 =>	x"06060606",
		1268 =>	x"06060606",
		1269 =>	x"06060606",
		1270 =>	x"06060606",
		1271 =>	x"06060606",
		1272 =>	x"06060606",
		1273 =>	x"06060606",
		1274 =>	x"06060606",
		1275 =>	x"06060606",
		1276 =>	x"06060606",
		1277 =>	x"06060606",
		1278 =>	x"06060606",
		1279 =>	x"06060606", -- IMG_16x16_bg51
		1280 =>	x"06060606",
		1281 =>	x"06060606",
		1282 =>	x"06060606",
		1283 =>	x"06060606",
		1284 =>	x"06060606",
		1285 =>	x"06060606",
		1286 =>	x"06060606",
		1287 =>	x"06060606",
		1288 =>	x"06060606",
		1289 =>	x"06060606",
		1290 =>	x"06060606",
		1291 =>	x"06060606",
		1292 =>	x"06060606",
		1293 =>	x"06060606",
		1294 =>	x"06060606",
		1295 =>	x"06060606",
		1296 =>	x"06060606",
		1297 =>	x"06060606",
		1298 =>	x"06060606",
		1299 =>	x"06060606",
		1300 =>	x"06060606",
		1301 =>	x"06060606",
		1302 =>	x"06060606",
		1303 =>	x"06060606",
		1304 =>	x"06060606",
		1305 =>	x"06060606",
		1306 =>	x"06060606",
		1307 =>	x"06060606",
		1308 =>	x"06060606",
		1309 =>	x"06060606",
		1310 =>	x"06060606",
		1311 =>	x"06060606",
		1312 =>	x"06060707",
		1313 =>	x"06060606",
		1314 =>	x"06060606",
		1315 =>	x"06060606",
		1316 =>	x"06060706",
		1317 =>	x"06060606",
		1318 =>	x"06060606",
		1319 =>	x"06060606",
		1320 =>	x"06060606",
		1321 =>	x"06060606",
		1322 =>	x"06060606",
		1323 =>	x"06060606",
		1324 =>	x"06060606",
		1325 =>	x"06060606",
		1326 =>	x"06060606",
		1327 =>	x"06060606",
		1328 =>	x"06060606",
		1329 =>	x"06060606",
		1330 =>	x"06060606",
		1331 =>	x"06060606",
		1332 =>	x"06060606",
		1333 =>	x"06060606",
		1334 =>	x"06060606",
		1335 =>	x"06060606",
		1336 =>	x"06060606",
		1337 =>	x"06060606",
		1338 =>	x"06060606",
		1339 =>	x"06060606",
		1340 =>	x"06060606",
		1341 =>	x"06060606",
		1342 =>	x"06060606",
		1343 =>	x"06060606", -- IMG_16x16_bg52
		1344 =>	x"06060606",
		1345 =>	x"06060606",
		1346 =>	x"06060606",
		1347 =>	x"06060606",
		1348 =>	x"06060606",
		1349 =>	x"06060606",
		1350 =>	x"06060606",
		1351 =>	x"06060606",
		1352 =>	x"06060606",
		1353 =>	x"06060606",
		1354 =>	x"06060607",
		1355 =>	x"06060606",
		1356 =>	x"06060606",
		1357 =>	x"06060606",
		1358 =>	x"06060607",
		1359 =>	x"06060606",
		1360 =>	x"06060606",
		1361 =>	x"06060606",
		1362 =>	x"06060606",
		1363 =>	x"06060606",
		1364 =>	x"06060606",
		1365 =>	x"06060606",
		1366 =>	x"06060606",
		1367 =>	x"06060606",
		1368 =>	x"06060606",
		1369 =>	x"06060606",
		1370 =>	x"06060606",
		1371 =>	x"06060606",
		1372 =>	x"06060606",
		1373 =>	x"06060606",
		1374 =>	x"06060606",
		1375 =>	x"06060606",
		1376 =>	x"06060606",
		1377 =>	x"06060606",
		1378 =>	x"06060606",
		1379 =>	x"06060606",
		1380 =>	x"06060606",
		1381 =>	x"06060606",
		1382 =>	x"06060606",
		1383 =>	x"06060606",
		1384 =>	x"06060606",
		1385 =>	x"06060606",
		1386 =>	x"06060606",
		1387 =>	x"06060606",
		1388 =>	x"06060606",
		1389 =>	x"06060606",
		1390 =>	x"06060606",
		1391 =>	x"06060606",
		1392 =>	x"06060606",
		1393 =>	x"06060606",
		1394 =>	x"06060606",
		1395 =>	x"06060606",
		1396 =>	x"06060606",
		1397 =>	x"06060606",
		1398 =>	x"06060606",
		1399 =>	x"06060606",
		1400 =>	x"06060606",
		1401 =>	x"06060606",
		1402 =>	x"06060606",
		1403 =>	x"06060606",
		1404 =>	x"06060606",
		1405 =>	x"06060606",
		1406 =>	x"06060606",
		1407 =>	x"00000000", -- IMG_16x16_black
		1408 =>	x"00000000",
		1409 =>	x"00000000",
		1410 =>	x"00000000",
		1411 =>	x"00000000",
		1412 =>	x"00000000",
		1413 =>	x"00000000",
		1414 =>	x"00000000",
		1415 =>	x"00000000",
		1416 =>	x"00000000",
		1417 =>	x"00000000",
		1418 =>	x"00000000",
		1419 =>	x"00000000",
		1420 =>	x"00000000",
		1421 =>	x"00000000",
		1422 =>	x"00000000",
		1423 =>	x"00000000",
		1424 =>	x"00000000",
		1425 =>	x"00000000",
		1426 =>	x"00000000",
		1427 =>	x"00000000",
		1428 =>	x"00000000",
		1429 =>	x"00000000",
		1430 =>	x"00000000",
		1431 =>	x"00000000",
		1432 =>	x"00000000",
		1433 =>	x"00000000",
		1434 =>	x"00000000",
		1435 =>	x"00000000",
		1436 =>	x"00000000",
		1437 =>	x"00000000",
		1438 =>	x"00000000",
		1439 =>	x"00000000",
		1440 =>	x"00000000",
		1441 =>	x"00000000",
		1442 =>	x"00000000",
		1443 =>	x"00000000",
		1444 =>	x"00000000",
		1445 =>	x"00000000",
		1446 =>	x"00000000",
		1447 =>	x"00000000",
		1448 =>	x"00000000",
		1449 =>	x"00000000",
		1450 =>	x"00000000",
		1451 =>	x"00000000",
		1452 =>	x"00000000",
		1453 =>	x"00000000",
		1454 =>	x"00000000",
		1455 =>	x"00000000",
		1456 =>	x"00000000",
		1457 =>	x"00000000",
		1458 =>	x"00000000",
		1459 =>	x"00000000",
		1460 =>	x"00000000",
		1461 =>	x"00000000",
		1462 =>	x"00000000",
		1463 =>	x"00000000",
		1464 =>	x"00000000",
		1465 =>	x"00000000",
		1466 =>	x"00000000",
		1467 =>	x"00000000",
		1468 =>	x"00000000",
		1469 =>	x"00000000",
		1470 =>	x"00000000",
		1471 =>	x"00000000", -- IMG_16x16_cursor
		1472 =>	x"00000000",
		1473 =>	x"00000000",
		1474 =>	x"00000000",
		1475 =>	x"00000000",
		1476 =>	x"00000008",
		1477 =>	x"00000000",
		1478 =>	x"00000000",
		1479 =>	x"00000000",
		1480 =>	x"00080808",
		1481 =>	x"08080000",
		1482 =>	x"00000000",
		1483 =>	x"00000008",
		1484 =>	x"08080808",
		1485 =>	x"08080808",
		1486 =>	x"00000000",
		1487 =>	x"00000808",
		1488 =>	x"08000008",
		1489 =>	x"00000808",
		1490 =>	x"08000000",
		1491 =>	x"00000808",
		1492 =>	x"00000008",
		1493 =>	x"00000008",
		1494 =>	x"08000000",
		1495 =>	x"00080800",
		1496 =>	x"00000008",
		1497 =>	x"00000000",
		1498 =>	x"08080000",
		1499 =>	x"00080800",
		1500 =>	x"00000008",
		1501 =>	x"00000000",
		1502 =>	x"08080000",
		1503 =>	x"08080809",
		1504 =>	x"0A080808",
		1505 =>	x"08080808",
		1506 =>	x"0A080800",
		1507 =>	x"00080800",
		1508 =>	x"00000008",
		1509 =>	x"00000000",
		1510 =>	x"08080000",
		1511 =>	x"00080800",
		1512 =>	x"00000008",
		1513 =>	x"00000000",
		1514 =>	x"08080000",
		1515 =>	x"00000808",
		1516 =>	x"00000008",
		1517 =>	x"00000008",
		1518 =>	x"08000000",
		1519 =>	x"00000808",
		1520 =>	x"08000008",
		1521 =>	x"00000808",
		1522 =>	x"08000000",
		1523 =>	x"00000008",
		1524 =>	x"08080808",
		1525 =>	x"08080808",
		1526 =>	x"00000000",
		1527 =>	x"00000000",
		1528 =>	x"00080808",
		1529 =>	x"08080000",
		1530 =>	x"00000000",
		1531 =>	x"00000000",
		1532 =>	x"00000008",
		1533 =>	x"00000000",
		1534 =>	x"00000000",
		1535 =>	x"00000000", -- IMG_16x16_four
		1536 =>	x"00000000",
		1537 =>	x"00000000",
		1538 =>	x"00000000",
		1539 =>	x"00000000",
		1540 =>	x"00000000",
		1541 =>	x"00000000",
		1542 =>	x"00000000",
		1543 =>	x"00000000",
		1544 =>	x"00000000",
		1545 =>	x"00000300",
		1546 =>	x"00000000",
		1547 =>	x"00000000",
		1548 =>	x"00000000",
		1549 =>	x"00030300",
		1550 =>	x"00000000",
		1551 =>	x"00000000",
		1552 =>	x"00000000",
		1553 =>	x"03000300",
		1554 =>	x"00000000",
		1555 =>	x"00000000",
		1556 =>	x"00000003",
		1557 =>	x"00000300",
		1558 =>	x"00000000",
		1559 =>	x"00000000",
		1560 =>	x"00000300",
		1561 =>	x"00000300",
		1562 =>	x"00000000",
		1563 =>	x"00000000",
		1564 =>	x"00030000",
		1565 =>	x"00000300",
		1566 =>	x"00000000",
		1567 =>	x"00000000",
		1568 =>	x"03030303",
		1569 =>	x"03030303",
		1570 =>	x"03000000",
		1571 =>	x"00000000",
		1572 =>	x"00000000",
		1573 =>	x"00000300",
		1574 =>	x"00000000",
		1575 =>	x"00000000",
		1576 =>	x"00000000",
		1577 =>	x"00000300",
		1578 =>	x"00000000",
		1579 =>	x"00000000",
		1580 =>	x"00000000",
		1581 =>	x"00000300",
		1582 =>	x"00000000",
		1583 =>	x"00000000",
		1584 =>	x"00000000",
		1585 =>	x"00000300",
		1586 =>	x"00000000",
		1587 =>	x"00000000",
		1588 =>	x"00000000",
		1589 =>	x"00000300",
		1590 =>	x"00000000",
		1591 =>	x"00000000",
		1592 =>	x"00000000",
		1593 =>	x"00000000",
		1594 =>	x"00000000",
		1595 =>	x"00000000",
		1596 =>	x"00000000",
		1597 =>	x"00000000",
		1598 =>	x"00000000",
		1599 =>	x"00000000", -- IMG_16x16_one
		1600 =>	x"00000000",
		1601 =>	x"00000000",
		1602 =>	x"00000000",
		1603 =>	x"00000000",
		1604 =>	x"00000000",
		1605 =>	x"00000000",
		1606 =>	x"00000000",
		1607 =>	x"00000000",
		1608 =>	x"00000000",
		1609 =>	x"03000000",
		1610 =>	x"00000000",
		1611 =>	x"00000000",
		1612 =>	x"00000003",
		1613 =>	x"03000000",
		1614 =>	x"00000000",
		1615 =>	x"00000000",
		1616 =>	x"00000300",
		1617 =>	x"03000000",
		1618 =>	x"00000000",
		1619 =>	x"00000000",
		1620 =>	x"00030000",
		1621 =>	x"03000000",
		1622 =>	x"00000000",
		1623 =>	x"00000000",
		1624 =>	x"03000000",
		1625 =>	x"03000000",
		1626 =>	x"00000000",
		1627 =>	x"00000000",
		1628 =>	x"00000000",
		1629 =>	x"03000000",
		1630 =>	x"00000000",
		1631 =>	x"00000000",
		1632 =>	x"00000000",
		1633 =>	x"03000000",
		1634 =>	x"00000000",
		1635 =>	x"00000000",
		1636 =>	x"00000000",
		1637 =>	x"03000000",
		1638 =>	x"00000000",
		1639 =>	x"00000000",
		1640 =>	x"00000000",
		1641 =>	x"03000000",
		1642 =>	x"00000000",
		1643 =>	x"00000000",
		1644 =>	x"00000000",
		1645 =>	x"03000000",
		1646 =>	x"00000000",
		1647 =>	x"00000000",
		1648 =>	x"00000000",
		1649 =>	x"03000000",
		1650 =>	x"00000000",
		1651 =>	x"00000000",
		1652 =>	x"00000000",
		1653 =>	x"00000000",
		1654 =>	x"00000000",
		1655 =>	x"00000000",
		1656 =>	x"00000000",
		1657 =>	x"00000000",
		1658 =>	x"00000000",
		1659 =>	x"00000000",
		1660 =>	x"00000000",
		1661 =>	x"00000000",
		1662 =>	x"00000000",
		1663 =>	x"00000000", -- IMG_16x16_pl00
		1664 =>	x"00000000",
		1665 =>	x"00000000",
		1666 =>	x"00000000",
		1667 =>	x"00000000",
		1668 =>	x"00000000",
		1669 =>	x"00000000",
		1670 =>	x"00000000",
		1671 =>	x"00000000",
		1672 =>	x"00000000",
		1673 =>	x"000B0000",
		1674 =>	x"00000000",
		1675 =>	x"00000000",
		1676 =>	x"00000000",
		1677 =>	x"0C0D0C00",
		1678 =>	x"00000000",
		1679 =>	x"00000000",
		1680 =>	x"0E0E000C",
		1681 =>	x"0303030C",
		1682 =>	x"0C000000",
		1683 =>	x"00000000",
		1684 =>	x"0E0E0E0C",
		1685 =>	x"0300030C",
		1686 =>	x"0C000000",
		1687 =>	x"00000000",
		1688 =>	x"000E0E0C",
		1689 =>	x"0303030C",
		1690 =>	x"0C000000",
		1691 =>	x"00000000",
		1692 =>	x"00000E0C",
		1693 =>	x"0C030C0C",
		1694 =>	x"0C000000",
		1695 =>	x"00000000",
		1696 =>	x"0000000C",
		1697 =>	x"0C0C0C0C",
		1698 =>	x"0C0C0000",
		1699 =>	x"00000000",
		1700 =>	x"00000000",
		1701 =>	x"0C0C0C0C",
		1702 =>	x"0C0C0C00",
		1703 =>	x"00000000",
		1704 =>	x"00000000",
		1705 =>	x"000C0C0C",
		1706 =>	x"0C0C0C00",
		1707 =>	x"00000000",
		1708 =>	x"00000000",
		1709 =>	x"000C0C00",
		1710 =>	x"00000000",
		1711 =>	x"00000000",
		1712 =>	x"00000000",
		1713 =>	x"00000008",
		1714 =>	x"08080808",
		1715 =>	x"00000000",
		1716 =>	x"00000000",
		1717 =>	x"00000808",
		1718 =>	x"08080808",
		1719 =>	x"00000000",
		1720 =>	x"00000000",
		1721 =>	x"00000808",
		1722 =>	x"08080808",
		1723 =>	x"00000000",
		1724 =>	x"00000808",
		1725 =>	x"08080808",
		1726 =>	x"08080808",
		1727 =>	x"00000000", -- IMG_16x16_pl01
		1728 =>	x"00000000",
		1729 =>	x"00000000",
		1730 =>	x"00000000",
		1731 =>	x"00000000",
		1732 =>	x"00000000",
		1733 =>	x"00000000",
		1734 =>	x"00000000",
		1735 =>	x"00000000",
		1736 =>	x"00000000",
		1737 =>	x"00000000",
		1738 =>	x"00000000",
		1739 =>	x"00000000",
		1740 =>	x"00000000",
		1741 =>	x"00000000",
		1742 =>	x"00000000",
		1743 =>	x"00000000",
		1744 =>	x"00000000",
		1745 =>	x"00000000",
		1746 =>	x"00000000",
		1747 =>	x"00000000",
		1748 =>	x"00000000",
		1749 =>	x"00000000",
		1750 =>	x"00000000",
		1751 =>	x"00000000",
		1752 =>	x"00000000",
		1753 =>	x"00000000",
		1754 =>	x"00000000",
		1755 =>	x"00000000",
		1756 =>	x"00000000",
		1757 =>	x"00000000",
		1758 =>	x"00000000",
		1759 =>	x"00000000",
		1760 =>	x"00000000",
		1761 =>	x"00000000",
		1762 =>	x"00000000",
		1763 =>	x"00000000",
		1764 =>	x"00000000",
		1765 =>	x"00000000",
		1766 =>	x"00000000",
		1767 =>	x"00000000",
		1768 =>	x"00000000",
		1769 =>	x"00000000",
		1770 =>	x"00000000",
		1771 =>	x"00000000",
		1772 =>	x"00000000",
		1773 =>	x"00000000",
		1774 =>	x"00000000",
		1775 =>	x"00000000",
		1776 =>	x"00000008",
		1777 =>	x"08000000",
		1778 =>	x"00000000",
		1779 =>	x"08000000",
		1780 =>	x"08080808",
		1781 =>	x"08080808",
		1782 =>	x"00000000",
		1783 =>	x"08080808",
		1784 =>	x"08080808",
		1785 =>	x"08080808",
		1786 =>	x"00000000",
		1787 =>	x"08080808",
		1788 =>	x"08080808",
		1789 =>	x"08080000",
		1790 =>	x"00000000",
		1791 =>	x"00000000", -- IMG_16x16_pl10
		1792 =>	x"08080808",
		1793 =>	x"08080808",
		1794 =>	x"08080808",
		1795 =>	x"00000008",
		1796 =>	x"08080808",
		1797 =>	x"08080808",
		1798 =>	x"08080808",
		1799 =>	x"00000808",
		1800 =>	x"08080808",
		1801 =>	x"08080808",
		1802 =>	x"08080808",
		1803 =>	x"00080808",
		1804 =>	x"08080808",
		1805 =>	x"08080808",
		1806 =>	x"08080808",
		1807 =>	x"00000808",
		1808 =>	x"08080808",
		1809 =>	x"08080808",
		1810 =>	x"08080808",
		1811 =>	x"00000008",
		1812 =>	x"08000808",
		1813 =>	x"00080808",
		1814 =>	x"08080808",
		1815 =>	x"00000000",
		1816 =>	x"00000000",
		1817 =>	x"00000000",
		1818 =>	x"08080808",
		1819 =>	x"00000000",
		1820 =>	x"00000000",
		1821 =>	x"00000000",
		1822 =>	x"00080808",
		1823 =>	x"00000000",
		1824 =>	x"00000000",
		1825 =>	x"00000000",
		1826 =>	x"00000808",
		1827 =>	x"00000000",
		1828 =>	x"00000000",
		1829 =>	x"00000000",
		1830 =>	x"00000000",
		1831 =>	x"00000000",
		1832 =>	x"00000000",
		1833 =>	x"00000000",
		1834 =>	x"00000000",
		1835 =>	x"00000000",
		1836 =>	x"00000000",
		1837 =>	x"00000000",
		1838 =>	x"00000000",
		1839 =>	x"00000000",
		1840 =>	x"00000000",
		1841 =>	x"00000000",
		1842 =>	x"00000000",
		1843 =>	x"00000000",
		1844 =>	x"00000000",
		1845 =>	x"00000000",
		1846 =>	x"00000000",
		1847 =>	x"00000000",
		1848 =>	x"00000000",
		1849 =>	x"00000000",
		1850 =>	x"00000000",
		1851 =>	x"00000000",
		1852 =>	x"00000000",
		1853 =>	x"00000000",
		1854 =>	x"00000000",
		1855 =>	x"08080808", -- IMG_16x16_pl11
		1856 =>	x"08080808",
		1857 =>	x"08080000",
		1858 =>	x"00000000",
		1859 =>	x"08080808",
		1860 =>	x"08080808",
		1861 =>	x"08000000",
		1862 =>	x"00000000",
		1863 =>	x"08080808",
		1864 =>	x"08080808",
		1865 =>	x"08000000",
		1866 =>	x"00000000",
		1867 =>	x"08080808",
		1868 =>	x"08080808",
		1869 =>	x"08000000",
		1870 =>	x"00000000",
		1871 =>	x"08080808",
		1872 =>	x"08080808",
		1873 =>	x"08080000",
		1874 =>	x"00000000",
		1875 =>	x"08080808",
		1876 =>	x"08080808",
		1877 =>	x"08080800",
		1878 =>	x"00000000",
		1879 =>	x"08080808",
		1880 =>	x"08080808",
		1881 =>	x"08080800",
		1882 =>	x"00000000",
		1883 =>	x"08080808",
		1884 =>	x"08080808",
		1885 =>	x"08080800",
		1886 =>	x"00000000",
		1887 =>	x"08080808",
		1888 =>	x"08080808",
		1889 =>	x"08000000",
		1890 =>	x"00000000",
		1891 =>	x"00000808",
		1892 =>	x"08000000",
		1893 =>	x"00000000",
		1894 =>	x"00000000",
		1895 =>	x"00000000",
		1896 =>	x"00000000",
		1897 =>	x"00000000",
		1898 =>	x"00000000",
		1899 =>	x"00000000",
		1900 =>	x"0000000E",
		1901 =>	x"0E000000",
		1902 =>	x"00000000",
		1903 =>	x"0000000E",
		1904 =>	x"0E00000E",
		1905 =>	x"0E0E0000",
		1906 =>	x"00000000",
		1907 =>	x"0000000E",
		1908 =>	x"0E0E0000",
		1909 =>	x"0E000000",
		1910 =>	x"00000000",
		1911 =>	x"00000000",
		1912 =>	x"0E0E0E00",
		1913 =>	x"00000000",
		1914 =>	x"00000000",
		1915 =>	x"00000000",
		1916 =>	x"000E0000",
		1917 =>	x"00000000",
		1918 =>	x"00000000",
		1919 =>	x"00000000", -- IMG_16x16_pr00
		1920 =>	x"00000000",
		1921 =>	x"00000000",
		1922 =>	x"00000000",
		1923 =>	x"00000000",
		1924 =>	x"00000000",
		1925 =>	x"00000000",
		1926 =>	x"00000000",
		1927 =>	x"00000000",
		1928 =>	x"00000000",
		1929 =>	x"00000000",
		1930 =>	x"0000000C",
		1931 =>	x"00000000",
		1932 =>	x"00000000",
		1933 =>	x"00000000",
		1934 =>	x"00000C0C",
		1935 =>	x"00000000",
		1936 =>	x"00000000",
		1937 =>	x"00000000",
		1938 =>	x"000C0C0C",
		1939 =>	x"00000000",
		1940 =>	x"00000000",
		1941 =>	x"00000000",
		1942 =>	x"000C0C0C",
		1943 =>	x"00000000",
		1944 =>	x"00000000",
		1945 =>	x"00000000",
		1946 =>	x"000C0C0C",
		1947 =>	x"00000000",
		1948 =>	x"00000000",
		1949 =>	x"00000000",
		1950 =>	x"0C0C0C0C",
		1951 =>	x"00000000",
		1952 =>	x"00000000",
		1953 =>	x"00000000",
		1954 =>	x"0C0C0C0C",
		1955 =>	x"00000000",
		1956 =>	x"00000000",
		1957 =>	x"00000000",
		1958 =>	x"000C0C0C",
		1959 =>	x"00000000",
		1960 =>	x"00000000",
		1961 =>	x"00000000",
		1962 =>	x"000C0C0C",
		1963 =>	x"00000000",
		1964 =>	x"00000000",
		1965 =>	x"00000000",
		1966 =>	x"00000000",
		1967 =>	x"00000000",
		1968 =>	x"00000000",
		1969 =>	x"00000000",
		1970 =>	x"00080808",
		1971 =>	x"00000000",
		1972 =>	x"00080808",
		1973 =>	x"00000000",
		1974 =>	x"08080808",
		1975 =>	x"00080808",
		1976 =>	x"08080808",
		1977 =>	x"08080808",
		1978 =>	x"08080808",
		1979 =>	x"00000808",
		1980 =>	x"08080808",
		1981 =>	x"08080808",
		1982 =>	x"08080808",
		1983 =>	x"00000000", -- IMG_16x16_pr01
		1984 =>	x"00000000",
		1985 =>	x"00000000",
		1986 =>	x"00000000",
		1987 =>	x"00000000",
		1988 =>	x"00000000",
		1989 =>	x"00000000",
		1990 =>	x"00000000",
		1991 =>	x"0C0C0000",
		1992 =>	x"00000000",
		1993 =>	x"00000000",
		1994 =>	x"00000000",
		1995 =>	x"0C030C0C",
		1996 =>	x"00000F0F",
		1997 =>	x"00000000",
		1998 =>	x"00000000",
		1999 =>	x"0303030C",
		2000 =>	x"0C0F0F0F",
		2001 =>	x"00000000",
		2002 =>	x"00000000",
		2003 =>	x"0300030C",
		2004 =>	x"0C0F0F0F",
		2005 =>	x"00000000",
		2006 =>	x"00000000",
		2007 =>	x"0303030C",
		2008 =>	x"0C0F0F00",
		2009 =>	x"00000000",
		2010 =>	x"00000000",
		2011 =>	x"0C030C0C",
		2012 =>	x"0C0F0000",
		2013 =>	x"00000000",
		2014 =>	x"00000000",
		2015 =>	x"0C0C0C0C",
		2016 =>	x"0C000000",
		2017 =>	x"00000000",
		2018 =>	x"00000000",
		2019 =>	x"0C0C0C0C",
		2020 =>	x"0C000000",
		2021 =>	x"00000000",
		2022 =>	x"00000000",
		2023 =>	x"0C0C0C0C",
		2024 =>	x"00000000",
		2025 =>	x"00000000",
		2026 =>	x"00000000",
		2027 =>	x"00000C00",
		2028 =>	x"00000000",
		2029 =>	x"00000000",
		2030 =>	x"00000000",
		2031 =>	x"08000000",
		2032 =>	x"00000000",
		2033 =>	x"00000000",
		2034 =>	x"00000000",
		2035 =>	x"08080800",
		2036 =>	x"00000000",
		2037 =>	x"00000000",
		2038 =>	x"00000000",
		2039 =>	x"08080808",
		2040 =>	x"00000000",
		2041 =>	x"00000000",
		2042 =>	x"00000000",
		2043 =>	x"08080808",
		2044 =>	x"08080808",
		2045 =>	x"00000000",
		2046 =>	x"00000000",
		2047 =>	x"00000808", -- IMG_16x16_pr10
		2048 =>	x"08080808",
		2049 =>	x"08080808",
		2050 =>	x"08080808",
		2051 =>	x"00000008",
		2052 =>	x"08080808",
		2053 =>	x"08080808",
		2054 =>	x"08080808",
		2055 =>	x"00000008",
		2056 =>	x"08080808",
		2057 =>	x"08080808",
		2058 =>	x"08080808",
		2059 =>	x"00000000",
		2060 =>	x"00080808",
		2061 =>	x"08080808",
		2062 =>	x"08080808",
		2063 =>	x"00000000",
		2064 =>	x"00000808",
		2065 =>	x"08080808",
		2066 =>	x"08080808",
		2067 =>	x"00000000",
		2068 =>	x"00000008",
		2069 =>	x"08080808",
		2070 =>	x"08080808",
		2071 =>	x"00000000",
		2072 =>	x"00000008",
		2073 =>	x"08080808",
		2074 =>	x"08080808",
		2075 =>	x"00000000",
		2076 =>	x"00000808",
		2077 =>	x"08080808",
		2078 =>	x"08080808",
		2079 =>	x"00000000",
		2080 =>	x"00000808",
		2081 =>	x"08080808",
		2082 =>	x"08080800",
		2083 =>	x"00000000",
		2084 =>	x"00080808",
		2085 =>	x"08080808",
		2086 =>	x"00000000",
		2087 =>	x"00000000",
		2088 =>	x"00000808",
		2089 =>	x"08080000",
		2090 =>	x"00000000",
		2091 =>	x"00000000",
		2092 =>	x"00000000",
		2093 =>	x"0000000E",
		2094 =>	x"0E000000",
		2095 =>	x"00000000",
		2096 =>	x"0000000E",
		2097 =>	x"0E000E0E",
		2098 =>	x"0E000000",
		2099 =>	x"00000000",
		2100 =>	x"00000E0E",
		2101 =>	x"0E000E0E",
		2102 =>	x"0E000000",
		2103 =>	x"00000000",
		2104 =>	x"0000000E",
		2105 =>	x"0000000E",
		2106 =>	x"00000000",
		2107 =>	x"00000000",
		2108 =>	x"00000000",
		2109 =>	x"00000000",
		2110 =>	x"00000000",
		2111 =>	x"08080808", -- IMG_16x16_pr11
		2112 =>	x"08080808",
		2113 =>	x"08080000",
		2114 =>	x"00000000",
		2115 =>	x"08080808",
		2116 =>	x"08080808",
		2117 =>	x"08080800",
		2118 =>	x"00000000",
		2119 =>	x"08080808",
		2120 =>	x"08080808",
		2121 =>	x"08080808",
		2122 =>	x"08000000",
		2123 =>	x"08080808",
		2124 =>	x"08080808",
		2125 =>	x"08080808",
		2126 =>	x"08080000",
		2127 =>	x"08080808",
		2128 =>	x"08080808",
		2129 =>	x"08080808",
		2130 =>	x"08080800",
		2131 =>	x"08080808",
		2132 =>	x"08080808",
		2133 =>	x"08080808",
		2134 =>	x"00000000",
		2135 =>	x"08080800",
		2136 =>	x"00080808",
		2137 =>	x"08080000",
		2138 =>	x"00000000",
		2139 =>	x"08000000",
		2140 =>	x"00000008",
		2141 =>	x"00000000",
		2142 =>	x"00000000",
		2143 =>	x"00000000",
		2144 =>	x"00000000",
		2145 =>	x"00000000",
		2146 =>	x"00000000",
		2147 =>	x"00000000",
		2148 =>	x"00000000",
		2149 =>	x"00000000",
		2150 =>	x"00000000",
		2151 =>	x"00000000",
		2152 =>	x"00000000",
		2153 =>	x"00000000",
		2154 =>	x"00000000",
		2155 =>	x"00000000",
		2156 =>	x"00000000",
		2157 =>	x"00000000",
		2158 =>	x"00000000",
		2159 =>	x"00000000",
		2160 =>	x"00000000",
		2161 =>	x"00000000",
		2162 =>	x"00000000",
		2163 =>	x"00000000",
		2164 =>	x"00000000",
		2165 =>	x"00000000",
		2166 =>	x"00000000",
		2167 =>	x"00000000",
		2168 =>	x"00000000",
		2169 =>	x"00000000",
		2170 =>	x"00000000",
		2171 =>	x"00000000",
		2172 =>	x"00000000",
		2173 =>	x"00000000",
		2174 =>	x"00000000",
		2175 =>	x"10010101", -- IMG_16x16_sky
		2176 =>	x"01010101",
		2177 =>	x"01010101",
		2178 =>	x"01010101",
		2179 =>	x"01010101",
		2180 =>	x"01010101",
		2181 =>	x"01010101",
		2182 =>	x"01010101",
		2183 =>	x"01010101",
		2184 =>	x"01010101",
		2185 =>	x"01010101",
		2186 =>	x"01010101",
		2187 =>	x"01010101",
		2188 =>	x"01010101",
		2189 =>	x"01010101",
		2190 =>	x"01010101",
		2191 =>	x"01010101",
		2192 =>	x"01010101",
		2193 =>	x"01010101",
		2194 =>	x"01010101",
		2195 =>	x"01010101",
		2196 =>	x"01010101",
		2197 =>	x"01010101",
		2198 =>	x"01010101",
		2199 =>	x"01010101",
		2200 =>	x"01010101",
		2201 =>	x"01010101",
		2202 =>	x"01010101",
		2203 =>	x"01010101",
		2204 =>	x"01010101",
		2205 =>	x"01010101",
		2206 =>	x"01010101",
		2207 =>	x"01010101",
		2208 =>	x"01010101",
		2209 =>	x"01010101",
		2210 =>	x"01010101",
		2211 =>	x"01010101",
		2212 =>	x"01010101",
		2213 =>	x"01010101",
		2214 =>	x"01010101",
		2215 =>	x"01010101",
		2216 =>	x"01010101",
		2217 =>	x"01010101",
		2218 =>	x"01010101",
		2219 =>	x"01010101",
		2220 =>	x"01010101",
		2221 =>	x"01010101",
		2222 =>	x"01010101",
		2223 =>	x"01010101",
		2224 =>	x"01010101",
		2225 =>	x"01010101",
		2226 =>	x"01010101",
		2227 =>	x"01010101",
		2228 =>	x"01010101",
		2229 =>	x"01010101",
		2230 =>	x"01010101",
		2231 =>	x"01010101",
		2232 =>	x"01010101",
		2233 =>	x"01010101",
		2234 =>	x"01010101",
		2235 =>	x"01010101",
		2236 =>	x"01010101",
		2237 =>	x"01010101",
		2238 =>	x"01010101",
		2239 =>	x"00000000", -- IMG_16x16_three
		2240 =>	x"00000000",
		2241 =>	x"00000000",
		2242 =>	x"00000000",
		2243 =>	x"00000000",
		2244 =>	x"00000000",
		2245 =>	x"00000000",
		2246 =>	x"00000000",
		2247 =>	x"00000003",
		2248 =>	x"03030303",
		2249 =>	x"03030300",
		2250 =>	x"00000000",
		2251 =>	x"00000000",
		2252 =>	x"00000000",
		2253 =>	x"00000300",
		2254 =>	x"00000000",
		2255 =>	x"00000000",
		2256 =>	x"00000000",
		2257 =>	x"00000300",
		2258 =>	x"00000000",
		2259 =>	x"00000000",
		2260 =>	x"00000000",
		2261 =>	x"00000300",
		2262 =>	x"00000000",
		2263 =>	x"00000000",
		2264 =>	x"00000000",
		2265 =>	x"00000300",
		2266 =>	x"00000000",
		2267 =>	x"00000003",
		2268 =>	x"03030303",
		2269 =>	x"03030300",
		2270 =>	x"00000000",
		2271 =>	x"00000000",
		2272 =>	x"00000000",
		2273 =>	x"00000300",
		2274 =>	x"00000000",
		2275 =>	x"00000000",
		2276 =>	x"00000000",
		2277 =>	x"00000300",
		2278 =>	x"00000000",
		2279 =>	x"00000000",
		2280 =>	x"00000000",
		2281 =>	x"00000300",
		2282 =>	x"00000000",
		2283 =>	x"00000000",
		2284 =>	x"00000000",
		2285 =>	x"00000300",
		2286 =>	x"00000000",
		2287 =>	x"00000003",
		2288 =>	x"03030303",
		2289 =>	x"03030300",
		2290 =>	x"00000000",
		2291 =>	x"00000000",
		2292 =>	x"00000000",
		2293 =>	x"00000000",
		2294 =>	x"00000000",
		2295 =>	x"00000000",
		2296 =>	x"00000000",
		2297 =>	x"00000000",
		2298 =>	x"00000000",
		2299 =>	x"00000000",
		2300 =>	x"00000000",
		2301 =>	x"00000000",
		2302 =>	x"00000000",
		2303 =>	x"00000000", -- IMG_16x16_two
		2304 =>	x"00000000",
		2305 =>	x"00000000",
		2306 =>	x"00000000",
		2307 =>	x"00000000",
		2308 =>	x"00000000",
		2309 =>	x"00000000",
		2310 =>	x"00000000",
		2311 =>	x"00000003",
		2312 =>	x"03030303",
		2313 =>	x"03030300",
		2314 =>	x"00000000",
		2315 =>	x"00000000",
		2316 =>	x"00000000",
		2317 =>	x"00000300",
		2318 =>	x"00000000",
		2319 =>	x"00000000",
		2320 =>	x"00000000",
		2321 =>	x"00000300",
		2322 =>	x"00000000",
		2323 =>	x"00000000",
		2324 =>	x"00000000",
		2325 =>	x"00000300",
		2326 =>	x"00000000",
		2327 =>	x"00000003",
		2328 =>	x"03030303",
		2329 =>	x"03030300",
		2330 =>	x"00000000",
		2331 =>	x"00000003",
		2332 =>	x"00000000",
		2333 =>	x"00000000",
		2334 =>	x"00000000",
		2335 =>	x"00000003",
		2336 =>	x"00000000",
		2337 =>	x"00000000",
		2338 =>	x"00000000",
		2339 =>	x"00000003",
		2340 =>	x"00000000",
		2341 =>	x"00000000",
		2342 =>	x"00000000",
		2343 =>	x"00000003",
		2344 =>	x"00000000",
		2345 =>	x"00000000",
		2346 =>	x"00000000",
		2347 =>	x"00000003",
		2348 =>	x"00000000",
		2349 =>	x"00000000",
		2350 =>	x"00000000",
		2351 =>	x"00000003",
		2352 =>	x"03030303",
		2353 =>	x"03030300",
		2354 =>	x"00000000",
		2355 =>	x"00000000",
		2356 =>	x"00000000",
		2357 =>	x"00000000",
		2358 =>	x"00000011",
		2359 =>	x"00000000",
		2360 =>	x"00000000",
		2361 =>	x"00000000",
		2362 =>	x"00000000",
		2363 =>	x"00000000",
		2364 =>	x"00000000",
		2365 =>	x"00000000",
		2366 =>	x"00000000",
		2367 =>	x"03030303", -- IMG_16x16_white
		2368 =>	x"03030303",
		2369 =>	x"03030303",
		2370 =>	x"03030303",
		2371 =>	x"03030303",
		2372 =>	x"03030303",
		2373 =>	x"03030303",
		2374 =>	x"03030303",
		2375 =>	x"03030303",
		2376 =>	x"03030303",
		2377 =>	x"03030303",
		2378 =>	x"03030303",
		2379 =>	x"03030303",
		2380 =>	x"03030303",
		2381 =>	x"03030303",
		2382 =>	x"03030303",
		2383 =>	x"03030303",
		2384 =>	x"03030303",
		2385 =>	x"03030303",
		2386 =>	x"03030303",
		2387 =>	x"03030303",
		2388 =>	x"03030303",
		2389 =>	x"03030303",
		2390 =>	x"03030303",
		2391 =>	x"03030303",
		2392 =>	x"03030303",
		2393 =>	x"03030303",
		2394 =>	x"03030303",
		2395 =>	x"03030303",
		2396 =>	x"03030303",
		2397 =>	x"03030303",
		2398 =>	x"03030303",
		2399 =>	x"03030303",
		2400 =>	x"03030303",
		2401 =>	x"03030303",
		2402 =>	x"03030303",
		2403 =>	x"03030303",
		2404 =>	x"03030303",
		2405 =>	x"03030303",
		2406 =>	x"03030303",
		2407 =>	x"03030303",
		2408 =>	x"03030303",
		2409 =>	x"03030303",
		2410 =>	x"03030303",
		2411 =>	x"03030303",
		2412 =>	x"03030303",
		2413 =>	x"03030303",
		2414 =>	x"03030303",
		2415 =>	x"03030303",
		2416 =>	x"03030303",
		2417 =>	x"03030303",
		2418 =>	x"03030303",
		2419 =>	x"03030303",
		2420 =>	x"03030303",
		2421 =>	x"03030303",
		2422 =>	x"03030303",
		2423 =>	x"03030303",
		2424 =>	x"03030303",
		2425 =>	x"03030303",
		2426 =>	x"03030303",
		2427 =>	x"03030303",
		2428 =>	x"03030303",
		2429 =>	x"03030303",
		2430 =>	x"03030303",
		2431 =>	x"00000000", -- IMG_16x16_zero
		2432 =>	x"00000000",
		2433 =>	x"00000000",
		2434 =>	x"00001200",
		2435 =>	x"00000000",
		2436 =>	x"00000000",
		2437 =>	x"00000000",
		2438 =>	x"00000000",
		2439 =>	x"00000000",
		2440 =>	x"03030303",
		2441 =>	x"03030300",
		2442 =>	x"00000000",
		2443 =>	x"00000000",
		2444 =>	x"03000000",
		2445 =>	x"00000300",
		2446 =>	x"00000000",
		2447 =>	x"00000000",
		2448 =>	x"03000000",
		2449 =>	x"00000300",
		2450 =>	x"00000000",
		2451 =>	x"00000000",
		2452 =>	x"03000000",
		2453 =>	x"00000300",
		2454 =>	x"00000000",
		2455 =>	x"00000000",
		2456 =>	x"03000000",
		2457 =>	x"00000300",
		2458 =>	x"00000000",
		2459 =>	x"00000000",
		2460 =>	x"03000000",
		2461 =>	x"00000300",
		2462 =>	x"00000000",
		2463 =>	x"00000000",
		2464 =>	x"03000000",
		2465 =>	x"00000300",
		2466 =>	x"00000000",
		2467 =>	x"00000000",
		2468 =>	x"03000000",
		2469 =>	x"00000300",
		2470 =>	x"00000000",
		2471 =>	x"00000000",
		2472 =>	x"03000000",
		2473 =>	x"00000300",
		2474 =>	x"00000000",
		2475 =>	x"00000000",
		2476 =>	x"03000000",
		2477 =>	x"00000300",
		2478 =>	x"00000000",
		2479 =>	x"00000000",
		2480 =>	x"03000000",
		2481 =>	x"00000300",
		2482 =>	x"00000000",
		2483 =>	x"00000000",
		2484 =>	x"03030303",
		2485 =>	x"03030300",
		2486 =>	x"00000000",
		2487 =>	x"00000000",
		2488 =>	x"00000000",
		2489 =>	x"00000000",
		2490 =>	x"00000000",
		2491 =>	x"00000000",
		2492 =>	x"00000000",
		2493 =>	x"00000000",
		2494 =>	x"00000000",


--			***** MAP *****


		2495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		2999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3215 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3216 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3217 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3218 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3219 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3220 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3221 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3222 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3223 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3224 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3225 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3226 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3227 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3228 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3229 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3230 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3231 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3232 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3233 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3234 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3235 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3236 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3237 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3238 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3239 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3240 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3241 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3242 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3243 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3244 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3245 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3246 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3247 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3248 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3249 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3250 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3251 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3252 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3253 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3254 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3255 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3308 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3309 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3312 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3313 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3314 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3315 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3316 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3317 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3318 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3319 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3320 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3321 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3322 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3323 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3324 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3325 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3326 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3327 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3328 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3329 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3330 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3331 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3332 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3333 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3334 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3335 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3388 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3389 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3392 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3393 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3394 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3395 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3396 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3397 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3398 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3399 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3400 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3401 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3402 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3403 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3404 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3405 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3406 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3407 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3408 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3409 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3410 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3411 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3412 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3413 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3414 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3415 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3439 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3466 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3467 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3487 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3488 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3489 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3490 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3546 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3547 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3567 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3568 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3569 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3570 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3626 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3627 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3647 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3648 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3649 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3650 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3706 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3707 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3727 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3728 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3729 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3730 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3786 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3787 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3807 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3808 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3809 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3810 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3866 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3867 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3887 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3888 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3889 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3890 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3946 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3947 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3967 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3968 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3969 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3970 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		3971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		3999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4026 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4027 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4047 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4048 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4049 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4050 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4106 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4107 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4108 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4109 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4123 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4124 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4125 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4126 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4127 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4128 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4129 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4130 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4188 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4189 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		4190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4415 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4416 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4417 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4418 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4419 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4420 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4421 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4422 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4423 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4424 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4425 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4426 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4427 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4428 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4429 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4430 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4431 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4432 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4433 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4434 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4435 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4436 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4437 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4438 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4439 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4440 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4441 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4442 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4443 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4444 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4445 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4446 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4447 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4448 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4449 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4450 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4451 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4452 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4453 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4454 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4455 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4495 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4496 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4497 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4498 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4499 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4500 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4501 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4502 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4503 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4504 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4505 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4506 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4507 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4508 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4509 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4510 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4511 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4512 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4513 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4514 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4515 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4516 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4517 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4518 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4519 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4520 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4521 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4522 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4523 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4524 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4525 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4526 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4527 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4528 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4529 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4530 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4531 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4532 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4533 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4534 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4535 =>	x"000000FF", -- z: 0 rot: 0 ptr: 255
		4536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		4999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5055 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		5056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5093 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		5094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5439 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		5440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5652 =>	x"0100023F", -- z: 1 rot: 0 ptr: 575
		5653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		5999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6295 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6296 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6297 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6298 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6299 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6300 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6301 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6302 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6303 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6304 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6305 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6306 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6307 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6308 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6309 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6310 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6311 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6312 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6313 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6314 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6315 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6316 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6317 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6318 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6319 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6320 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6321 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6322 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6323 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6324 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6325 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6326 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6327 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6328 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6329 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6330 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6331 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6332 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6333 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6334 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6335 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6336 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6337 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6338 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6339 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6340 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6341 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6342 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6343 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6344 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6345 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6346 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6347 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6348 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6349 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6350 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6351 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6352 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6353 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6354 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6355 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6356 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6357 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6358 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6359 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6360 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6361 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6362 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6363 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6364 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6365 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6366 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6367 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6368 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6369 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6370 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6371 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6372 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6373 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6374 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6375 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6376 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6377 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6378 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6379 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6380 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6381 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6382 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6383 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6384 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6385 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6386 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6387 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6388 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6389 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6390 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6391 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6392 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6393 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6394 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6395 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6396 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6397 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6398 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6399 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6400 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6401 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6402 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6403 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6404 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6405 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6406 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6407 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6408 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6409 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6410 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6411 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6412 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6413 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6414 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6415 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6416 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6417 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6418 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6419 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6420 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6421 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6422 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6423 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6424 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6425 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6426 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6427 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6428 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6429 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6430 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6431 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6432 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6433 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6434 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6435 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6436 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6437 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6438 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6439 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6440 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6441 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6442 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6443 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6444 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6445 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6446 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6447 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6448 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6449 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6450 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6451 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6452 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6453 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6454 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6455 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6456 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6457 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6458 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6459 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6460 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6461 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6462 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6463 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6464 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6465 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6466 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6467 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6468 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6469 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6470 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6471 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6472 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6473 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6474 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6475 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6476 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6477 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6478 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6479 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6480 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6481 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6482 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6483 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6484 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6485 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6486 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6487 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6488 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6489 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6490 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6491 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6492 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6493 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6494 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6495 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6496 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6497 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6498 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6499 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6500 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6501 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6502 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6503 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6504 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6505 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6506 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6507 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6508 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6509 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6510 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6511 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6512 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6513 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6514 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6515 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6516 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6517 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6518 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6519 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6520 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6521 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6522 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6523 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6524 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6525 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6526 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6527 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6528 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6529 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6530 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6531 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6532 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6533 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6534 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6535 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6536 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6537 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6538 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6539 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6540 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6541 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6542 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6543 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6544 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6545 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6546 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6547 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6548 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6549 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6550 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6551 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6552 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6553 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6554 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6555 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6556 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6557 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6558 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6559 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6560 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6561 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6562 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6563 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6564 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6565 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6566 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6567 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6568 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6569 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6570 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6571 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6572 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6573 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6574 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6575 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6576 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6577 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6578 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6579 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6580 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6581 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6582 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6583 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6584 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6585 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6586 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6587 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6588 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6589 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6590 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6591 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6592 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6593 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6594 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6595 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6596 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6597 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6598 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6599 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6600 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6601 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6602 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6603 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6604 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6605 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6606 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6607 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6608 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6609 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6610 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6611 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6612 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6613 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6614 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6615 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6616 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6617 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6618 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6619 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6620 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6621 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6622 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6623 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6624 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6625 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6626 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6627 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6628 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6629 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6630 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6631 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6632 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6633 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6634 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6635 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6636 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6637 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6638 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6639 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6640 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6641 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6642 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6643 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6644 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6645 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6646 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6647 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6648 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6649 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6650 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6651 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6652 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6653 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6654 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6655 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6656 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6657 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6658 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6659 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6660 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6661 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6662 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6663 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6664 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6665 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6666 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6667 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6668 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6669 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6670 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6671 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6672 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6673 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6674 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6675 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6676 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6677 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6678 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6679 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6680 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6681 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6682 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6683 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6684 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6685 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6686 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6687 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6688 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6689 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6690 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6691 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6692 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6693 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6694 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6695 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6696 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6697 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6698 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6699 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6700 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6701 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6702 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6703 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6704 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6705 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6706 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6707 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6708 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6709 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6710 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6711 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6712 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6713 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6714 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6715 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6716 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6717 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6718 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6719 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6720 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6721 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6722 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6723 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6724 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6725 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6726 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6727 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6728 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6729 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6730 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6731 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6732 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6733 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6734 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6735 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6736 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6737 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6738 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6739 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6740 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6741 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6742 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6743 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6744 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6745 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6746 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6747 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6748 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6749 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6750 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6751 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6752 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6753 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6754 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6755 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6756 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6757 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6758 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6759 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6760 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6761 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6762 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6763 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6764 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6765 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6766 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6767 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6768 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6769 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6770 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6771 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6772 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6773 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6774 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6775 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6776 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6777 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6778 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6779 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6780 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6781 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6782 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6783 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6784 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6785 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6786 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6787 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6788 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6789 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6790 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6791 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6792 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6793 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6794 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6795 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6796 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6797 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6798 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6799 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6800 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6801 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6802 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6803 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6804 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6805 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6806 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6807 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6808 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6809 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6810 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6811 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6812 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6813 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6814 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6815 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6816 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6817 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6818 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6819 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6820 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6821 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6822 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6823 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6824 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6825 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6826 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6827 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6828 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6829 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6830 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6831 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6832 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6833 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6834 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6835 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6836 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6837 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6838 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6839 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6840 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6841 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6842 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6843 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6844 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6845 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6846 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6847 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6848 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6849 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6850 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6851 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6852 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6853 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6854 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6855 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6856 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6857 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6858 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6859 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6860 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6861 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6862 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6863 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6864 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6865 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6866 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6867 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6868 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6869 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6870 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6871 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6872 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6873 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6874 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6875 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6876 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6877 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6878 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6879 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6880 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6881 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6882 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6883 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6884 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6885 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6886 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6887 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6888 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6889 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6890 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6891 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6892 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6893 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6894 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6895 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6896 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6897 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6898 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6899 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6900 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6901 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6902 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6903 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6904 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6905 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6906 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6907 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6908 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6909 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6910 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6911 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6912 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6913 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6914 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6915 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6916 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6917 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6918 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6919 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6920 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6921 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6922 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6923 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6924 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6925 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6926 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6927 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6928 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6929 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6930 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6931 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6932 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6933 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6934 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6935 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6936 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6937 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6938 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6939 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6940 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6941 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6942 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6943 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6944 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6945 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6946 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6947 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6948 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6949 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6950 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6951 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6952 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6953 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6954 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6955 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6956 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6957 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6958 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6959 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6960 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6961 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6962 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6963 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6964 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6965 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6966 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6967 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6968 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6969 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6970 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6971 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6972 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6973 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6974 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6975 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6976 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6977 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6978 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6979 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6980 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6981 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6982 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6983 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6984 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6985 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6986 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6987 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6988 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6989 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6990 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6991 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6992 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6993 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6994 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6995 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6996 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6997 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6998 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		6999 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7000 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7001 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7002 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7003 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7004 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7005 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7006 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7007 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7008 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7009 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7010 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7011 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7012 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7013 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7014 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7015 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7016 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7017 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7018 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7019 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7020 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7021 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7022 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7023 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7024 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7025 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7026 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7027 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7028 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7029 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7030 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7031 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7032 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7033 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7034 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7035 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7036 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7037 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7038 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7039 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7040 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7041 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7042 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7043 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7044 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7045 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7046 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7047 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7048 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7049 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7050 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7051 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7052 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7053 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7054 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7055 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7056 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7057 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7058 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7059 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7060 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7061 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7062 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7063 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7064 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7065 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7066 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7067 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7068 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7069 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7070 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7071 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7072 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7073 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7074 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7075 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7076 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7077 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7078 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7079 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7080 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7081 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7082 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7083 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7084 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7085 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7086 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7087 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7088 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7089 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7090 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7091 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7092 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7093 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7094 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7095 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7096 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7097 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7098 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7099 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7100 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7101 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7102 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7103 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7104 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7105 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7106 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7107 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7108 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7109 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7110 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7111 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7112 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7113 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7114 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7115 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7116 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7117 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7118 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7119 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7120 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7121 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7122 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7123 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7124 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7125 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7126 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7127 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7128 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7129 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7130 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7131 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7132 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7133 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7134 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7135 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7136 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7137 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7138 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7139 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7140 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7141 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7142 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7143 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7144 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7145 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7146 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7147 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7148 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7149 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7150 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7151 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7152 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7153 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7154 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7155 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7156 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7157 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7158 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7159 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7160 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7161 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7162 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7163 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7164 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7165 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7166 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7167 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7168 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7169 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7170 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7171 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7172 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7173 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7174 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7175 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7176 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7177 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7178 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7179 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7180 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7181 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7182 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7183 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7184 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7185 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7186 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7187 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7188 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7189 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7190 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7191 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7192 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7193 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7194 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7195 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7196 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7197 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7198 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7199 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7200 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7201 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7202 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7203 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7204 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7205 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7206 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7207 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7208 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7209 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7210 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7211 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7212 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7213 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7214 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7215 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7216 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7217 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7218 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7219 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7220 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7221 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7222 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7223 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7224 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7225 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7226 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7227 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7228 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7229 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7230 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7231 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7232 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7233 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7234 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7235 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7236 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7237 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7238 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7239 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7240 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7241 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7242 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7243 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7244 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7245 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7246 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7247 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7248 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7249 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7250 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7251 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7252 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7253 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7254 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7255 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7256 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7257 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7258 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7259 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7260 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7261 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7262 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7263 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7264 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7265 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7266 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7267 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7268 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7269 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7270 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7271 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7272 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7273 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7274 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7275 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7276 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7277 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7278 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7279 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7280 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7281 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7282 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7283 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7284 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7285 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7286 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7287 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7288 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7289 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7290 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7291 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7292 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7293 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		7294 =>	x"0000017F", -- z: 0 rot: 0 ptr: 383
		others => x"00000000"

	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;